LIBRARY IEEE;
LIBRARY WORK;
USE WORK.UTILS.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY datapath IS
	PORT(
		-- entradas
		clock, reset: IN  STD_LOGIC;
		data_in		: IN  STD_LOGIC_VECTOR(n_bits - 1 DOWNTO 0);
		c 				: IN  STD_LOGIC_VECTOR(28 DOWNTO 0);
		-- flags
		N,Z,Ov,Cout : OUT STD_LOGIC;
		
		-- saida dados
		data_out		: OUT STD_LOGIC_VECTOR(n_bits - 1 DOWNTO 0)
	
	);
END datapath;

ARCHITECTURE behavior OF datapath IS
	-- sinais para a saida dos muxs 2:1 que selecionam o dado de entrada para os registradores
	SIGNAL saidas_mux_2_1: matriz_8bits;
	
	-- sinal para a saida dos registradores, que são conectados aos mux 8:1
	SIGNAL saidas_regs: matriz_8bits;
	
	-- sinal para a saida dos muxs 8:1, que são conectados as ulas
	SIGNAL saidas_mux_8_1: matriz_8bits_2;
	
	-- sinal para a saida das ulas
	SIGNAL saida_ula_1, saida_ula_2: STD_LOGIC_VECTOR(n_bits - 1 DOWNTO 0);
	
BEGIN
	-- TESTE
	
	data_out <= saidas_mux_8_1(2);
	
	-- cria os mux 2 pra 1
	for_mux_2_1: FOR i IN 0 TO n_bits - 1 GENERATE
		muxes_2_1: mux_2_1 PORT MAP(
							in_0 => data_in, 
							in_1 => saida_ula_2, 
							sel => c(i), 
							saida => saidas_mux_2_1(i)
						);
	END GENERATE;
	
	
	-- cria os registradores de 8 bits
	for_regs: FOR i IN 0 TO n_bits - 1 GENERATE
		regs: registrador PORT MAP(
										data => saidas_mux_2_1(i),
										clock => clock,
										clear => reset,
										enable => c(8 + i),
										q => saidas_regs(i)
				);
	END GENERATE for_regs;
	
	--cria os mux de 8 para 1, conectados as portas das ulas
	for_mux_8_1: FOR i IN 0 TO 2 GENERATE
		muxs_8_1: mux_8_1 PORT MAP(
						in_0 => saidas_regs(0),
						in_1 => saidas_regs(1),
						in_2 => saidas_regs(2),
						in_3 => saidas_regs(3),
						in_4 => saidas_regs(4),
						in_5 => saidas_regs(5),
						in_6 => saidas_regs(6),
						in_7 => saidas_regs(7),
						sel => c((18 + (i * 3)) DOWNTO (16 + (i * 3))),
						saida => saidas_mux_8_1(i)
					);
	END GENERATE for_mux_8_1;
	
	primeira_ula: 
	ula1 PORT MAP (
		a => saidas_mux_8_1(1),
		b => saidas_mux_8_1(2),
		op => c(26 DOWNTO 25),
		Ov => Ov,
		Cout => Cout,
		saida => saida_ula_1
	);
	
	segunda_ula: 
	ula2 PORT MAP (
		c => saidas_mux_8_1(0),
		d => saida_ula_1,
		op => c(28 DOWNTO 27),
		N => N,
		Z => Z,
		saida => saida_ula_2
	);
	
END behavior;